/*
 * rom_sine_cosine_360x16.v
 */

module rom_sine_cosine_360x16 (
    input      [8:0]  angle,        // 9-bit angle input (0-359)
    output reg [15:0] sine_out,     // 16-bit output for sine
    output reg [15:0] cosine_out    // 16-bit output for cosine
);

  // ROM content in arrays for sine and cosine
  reg [15:0] sine_table [0:359];
  reg [15:0] cosine_table [0:359];

  initial begin
    sine_table[0] = 16'h0000;  // Angle 0°
    sine_table[1] = 16'h023B;  // Angle 1°
    sine_table[2] = 16'h0477;  // Angle 2°
    sine_table[3] = 16'h06B2;  // Angle 3°
    sine_table[4] = 16'h08ED;  // Angle 4°
    sine_table[5] = 16'h0B27;  // Angle 5°
    sine_table[6] = 16'h0D61;  // Angle 6°
    sine_table[7] = 16'h0F99;  // Angle 7°
    sine_table[8] = 16'h11D0;  // Angle 8°
    sine_table[9] = 16'h1406;  // Angle 9°
    sine_table[10] = 16'h163A;  // Angle 10°
    sine_table[11] = 16'h186C;  // Angle 11°
    sine_table[12] = 16'h1A9C;  // Angle 12°
    sine_table[13] = 16'h1CCB;  // Angle 13°
    sine_table[14] = 16'h1EF7;  // Angle 14°
    sine_table[15] = 16'h2120;  // Angle 15°
    sine_table[16] = 16'h2348;  // Angle 16°
    sine_table[17] = 16'h256C;  // Angle 17°
    sine_table[18] = 16'h278D;  // Angle 18°
    sine_table[19] = 16'h29AC;  // Angle 19°
    sine_table[20] = 16'h2BC7;  // Angle 20°
    sine_table[21] = 16'h2DDF;  // Angle 21°
    sine_table[22] = 16'h2FF3;  // Angle 22°
    sine_table[23] = 16'h3203;  // Angle 23°
    sine_table[24] = 16'h340F;  // Angle 24°
    sine_table[25] = 16'h3618;  // Angle 25°
    sine_table[26] = 16'h381C;  // Angle 26°
    sine_table[27] = 16'h3A1C;  // Angle 27°
    sine_table[28] = 16'h3C17;  // Angle 28°
    sine_table[29] = 16'h3E0E;  // Angle 29°
    sine_table[30] = 16'h3FFF;  // Angle 30°
    sine_table[31] = 16'h41EC;  // Angle 31°
    sine_table[32] = 16'h43D4;  // Angle 32°
    sine_table[33] = 16'h45B6;  // Angle 33°
    sine_table[34] = 16'h4793;  // Angle 34°
    sine_table[35] = 16'h496A;  // Angle 35°
    sine_table[36] = 16'h4B3C;  // Angle 36°
    sine_table[37] = 16'h4D08;  // Angle 37°
    sine_table[38] = 16'h4ECD;  // Angle 38°
    sine_table[39] = 16'h508D;  // Angle 39°
    sine_table[40] = 16'h5246;  // Angle 40°
    sine_table[41] = 16'h53F9;  // Angle 41°
    sine_table[42] = 16'h55A6;  // Angle 42°
    sine_table[43] = 16'h574B;  // Angle 43°
    sine_table[44] = 16'h58EA;  // Angle 44°
    sine_table[45] = 16'h5A82;  // Angle 45°
    sine_table[46] = 16'h5C13;  // Angle 46°
    sine_table[47] = 16'h5D9C;  // Angle 47°
    sine_table[48] = 16'h5F1F;  // Angle 48°
    sine_table[49] = 16'h609A;  // Angle 49°
    sine_table[50] = 16'h620D;  // Angle 50°
    sine_table[51] = 16'h6379;  // Angle 51°
    sine_table[52] = 16'h64DD;  // Angle 52°
    sine_table[53] = 16'h6639;  // Angle 53°
    sine_table[54] = 16'h678D;  // Angle 54°
    sine_table[55] = 16'h68D9;  // Angle 55°
    sine_table[56] = 16'h6A1D;  // Angle 56°
    sine_table[57] = 16'h6B59;  // Angle 57°
    sine_table[58] = 16'h6C8C;  // Angle 58°
    sine_table[59] = 16'h6DB7;  // Angle 59°
    sine_table[60] = 16'h6ED9;  // Angle 60°
    sine_table[61] = 16'h6FF3;  // Angle 61°
    sine_table[62] = 16'h7104;  // Angle 62°
    sine_table[63] = 16'h720C;  // Angle 63°
    sine_table[64] = 16'h730B;  // Angle 64°
    sine_table[65] = 16'h7401;  // Angle 65°
    sine_table[66] = 16'h74EF;  // Angle 66°
    sine_table[67] = 16'h75D3;  // Angle 67°
    sine_table[68] = 16'h76AD;  // Angle 68°
    sine_table[69] = 16'h777F;  // Angle 69°
    sine_table[70] = 16'h7847;  // Angle 70°
    sine_table[71] = 16'h7906;  // Angle 71°
    sine_table[72] = 16'h79BC;  // Angle 72°
    sine_table[73] = 16'h7A68;  // Angle 73°
    sine_table[74] = 16'h7B0A;  // Angle 74°
    sine_table[75] = 16'h7BA3;  // Angle 75°
    sine_table[76] = 16'h7C32;  // Angle 76°
    sine_table[77] = 16'h7CB8;  // Angle 77°
    sine_table[78] = 16'h7D33;  // Angle 78°
    sine_table[79] = 16'h7DA5;  // Angle 79°
    sine_table[80] = 16'h7E0E;  // Angle 80°
    sine_table[81] = 16'h7E6C;  // Angle 81°
    sine_table[82] = 16'h7EC1;  // Angle 82°
    sine_table[83] = 16'h7F0B;  // Angle 83°
    sine_table[84] = 16'h7F4C;  // Angle 84°
    sine_table[85] = 16'h7F83;  // Angle 85°
    sine_table[86] = 16'h7FB0;  // Angle 86°
    sine_table[87] = 16'h7FD3;  // Angle 87°
    sine_table[88] = 16'h7FEC;  // Angle 88°
    sine_table[89] = 16'h7FFB;  // Angle 89°
    sine_table[90] = 16'h7FFF;  // Angle 90°
    sine_table[91] = 16'h7FFB;  // Angle 91°
    sine_table[92] = 16'h7FEC;  // Angle 92°
    sine_table[93] = 16'h7FD3;  // Angle 93°
    sine_table[94] = 16'h7FB0;  // Angle 94°
    sine_table[95] = 16'h7F83;  // Angle 95°
    sine_table[96] = 16'h7F4C;  // Angle 96°
    sine_table[97] = 16'h7F0B;  // Angle 97°
    sine_table[98] = 16'h7EC1;  // Angle 98°
    sine_table[99] = 16'h7E6C;  // Angle 99°
    sine_table[100] = 16'h7E0E;  // Angle 100°
    sine_table[101] = 16'h7DA5;  // Angle 101°
    sine_table[102] = 16'h7D33;  // Angle 102°
    sine_table[103] = 16'h7CB8;  // Angle 103°
    sine_table[104] = 16'h7C32;  // Angle 104°
    sine_table[105] = 16'h7BA3;  // Angle 105°
    sine_table[106] = 16'h7B0A;  // Angle 106°
    sine_table[107] = 16'h7A68;  // Angle 107°
    sine_table[108] = 16'h79BC;  // Angle 108°
    sine_table[109] = 16'h7906;  // Angle 109°
    sine_table[110] = 16'h7847;  // Angle 110°
    sine_table[111] = 16'h777F;  // Angle 111°
    sine_table[112] = 16'h76AD;  // Angle 112°
    sine_table[113] = 16'h75D3;  // Angle 113°
    sine_table[114] = 16'h74EF;  // Angle 114°
    sine_table[115] = 16'h7401;  // Angle 115°
    sine_table[116] = 16'h730B;  // Angle 116°
    sine_table[117] = 16'h720C;  // Angle 117°
    sine_table[118] = 16'h7104;  // Angle 118°
    sine_table[119] = 16'h6FF3;  // Angle 119°
    sine_table[120] = 16'h6ED9;  // Angle 120°
    sine_table[121] = 16'h6DB7;  // Angle 121°
    sine_table[122] = 16'h6C8C;  // Angle 122°
    sine_table[123] = 16'h6B59;  // Angle 123°
    sine_table[124] = 16'h6A1D;  // Angle 124°
    sine_table[125] = 16'h68D9;  // Angle 125°
    sine_table[126] = 16'h678D;  // Angle 126°
    sine_table[127] = 16'h6639;  // Angle 127°
    sine_table[128] = 16'h64DD;  // Angle 128°
    sine_table[129] = 16'h6379;  // Angle 129°
    sine_table[130] = 16'h620D;  // Angle 130°
    sine_table[131] = 16'h609A;  // Angle 131°
    sine_table[132] = 16'h5F1F;  // Angle 132°
    sine_table[133] = 16'h5D9C;  // Angle 133°
    sine_table[134] = 16'h5C13;  // Angle 134°
    sine_table[135] = 16'h5A82;  // Angle 135°
    sine_table[136] = 16'h58EA;  // Angle 136°
    sine_table[137] = 16'h574B;  // Angle 137°
    sine_table[138] = 16'h55A6;  // Angle 138°
    sine_table[139] = 16'h53F9;  // Angle 139°
    sine_table[140] = 16'h5246;  // Angle 140°
    sine_table[141] = 16'h508D;  // Angle 141°
    sine_table[142] = 16'h4ECD;  // Angle 142°
    sine_table[143] = 16'h4D08;  // Angle 143°
    sine_table[144] = 16'h4B3C;  // Angle 144°
    sine_table[145] = 16'h496A;  // Angle 145°
    sine_table[146] = 16'h4793;  // Angle 146°
    sine_table[147] = 16'h45B6;  // Angle 147°
    sine_table[148] = 16'h43D4;  // Angle 148°
    sine_table[149] = 16'h41EC;  // Angle 149°
    sine_table[150] = 16'h3FFF;  // Angle 150°
    sine_table[151] = 16'h3E0E;  // Angle 151°
    sine_table[152] = 16'h3C17;  // Angle 152°
    sine_table[153] = 16'h3A1C;  // Angle 153°
    sine_table[154] = 16'h381C;  // Angle 154°
    sine_table[155] = 16'h3618;  // Angle 155°
    sine_table[156] = 16'h340F;  // Angle 156°
    sine_table[157] = 16'h3203;  // Angle 157°
    sine_table[158] = 16'h2FF3;  // Angle 158°
    sine_table[159] = 16'h2DDF;  // Angle 159°
    sine_table[160] = 16'h2BC7;  // Angle 160°
    sine_table[161] = 16'h29AC;  // Angle 161°
    sine_table[162] = 16'h278D;  // Angle 162°
    sine_table[163] = 16'h256C;  // Angle 163°
    sine_table[164] = 16'h2348;  // Angle 164°
    sine_table[165] = 16'h2120;  // Angle 165°
    sine_table[166] = 16'h1EF7;  // Angle 166°
    sine_table[167] = 16'h1CCB;  // Angle 167°
    sine_table[168] = 16'h1A9C;  // Angle 168°
    sine_table[169] = 16'h186C;  // Angle 169°
    sine_table[170] = 16'h163A;  // Angle 170°
    sine_table[171] = 16'h1406;  // Angle 171°
    sine_table[172] = 16'h11D0;  // Angle 172°
    sine_table[173] = 16'h0F99;  // Angle 173°
    sine_table[174] = 16'h0D61;  // Angle 174°
    sine_table[175] = 16'h0B27;  // Angle 175°
    sine_table[176] = 16'h08ED;  // Angle 176°
    sine_table[177] = 16'h06B2;  // Angle 177°
    sine_table[178] = 16'h0477;  // Angle 178°
    sine_table[179] = 16'h023B;  // Angle 179°
    sine_table[180] = 16'h0000;  // Angle 180°
    sine_table[181] = 16'hFDC5;  // Angle 181°
    sine_table[182] = 16'hFB89;  // Angle 182°
    sine_table[183] = 16'hF94E;  // Angle 183°
    sine_table[184] = 16'hF713;  // Angle 184°
    sine_table[185] = 16'hF4D9;  // Angle 185°
    sine_table[186] = 16'hF29F;  // Angle 186°
    sine_table[187] = 16'hF067;  // Angle 187°
    sine_table[188] = 16'hEE30;  // Angle 188°
    sine_table[189] = 16'hEBFA;  // Angle 189°
    sine_table[190] = 16'hE9C6;  // Angle 190°
    sine_table[191] = 16'hE794;  // Angle 191°
    sine_table[192] = 16'hE564;  // Angle 192°
    sine_table[193] = 16'hE335;  // Angle 193°
    sine_table[194] = 16'hE109;  // Angle 194°
    sine_table[195] = 16'hDEE0;  // Angle 195°
    sine_table[196] = 16'hDCB8;  // Angle 196°
    sine_table[197] = 16'hDA94;  // Angle 197°
    sine_table[198] = 16'hD873;  // Angle 198°
    sine_table[199] = 16'hD654;  // Angle 199°
    sine_table[200] = 16'hD439;  // Angle 200°
    sine_table[201] = 16'hD221;  // Angle 201°
    sine_table[202] = 16'hD00D;  // Angle 202°
    sine_table[203] = 16'hCDFD;  // Angle 203°
    sine_table[204] = 16'hCBF1;  // Angle 204°
    sine_table[205] = 16'hC9E8;  // Angle 205°
    sine_table[206] = 16'hC7E4;  // Angle 206°
    sine_table[207] = 16'hC5E4;  // Angle 207°
    sine_table[208] = 16'hC3E9;  // Angle 208°
    sine_table[209] = 16'hC1F2;  // Angle 209°
    sine_table[210] = 16'hC000;  // Angle 210°
    sine_table[211] = 16'hBE14;  // Angle 211°
    sine_table[212] = 16'hBC2C;  // Angle 212°
    sine_table[213] = 16'hBA4A;  // Angle 213°
    sine_table[214] = 16'hB86D;  // Angle 214°
    sine_table[215] = 16'hB696;  // Angle 215°
    sine_table[216] = 16'hB4C4;  // Angle 216°
    sine_table[217] = 16'hB2F8;  // Angle 217°
    sine_table[218] = 16'hB133;  // Angle 218°
    sine_table[219] = 16'hAF73;  // Angle 219°
    sine_table[220] = 16'hADBA;  // Angle 220°
    sine_table[221] = 16'hAC07;  // Angle 221°
    sine_table[222] = 16'hAA5A;  // Angle 222°
    sine_table[223] = 16'hA8B5;  // Angle 223°
    sine_table[224] = 16'hA716;  // Angle 224°
    sine_table[225] = 16'hA57E;  // Angle 225°
    sine_table[226] = 16'hA3ED;  // Angle 226°
    sine_table[227] = 16'hA264;  // Angle 227°
    sine_table[228] = 16'hA0E1;  // Angle 228°
    sine_table[229] = 16'h9F66;  // Angle 229°
    sine_table[230] = 16'h9DF3;  // Angle 230°
    sine_table[231] = 16'h9C87;  // Angle 231°
    sine_table[232] = 16'h9B23;  // Angle 232°
    sine_table[233] = 16'h99C7;  // Angle 233°
    sine_table[234] = 16'h9873;  // Angle 234°
    sine_table[235] = 16'h9727;  // Angle 235°
    sine_table[236] = 16'h95E3;  // Angle 236°
    sine_table[237] = 16'h94A7;  // Angle 237°
    sine_table[238] = 16'h9374;  // Angle 238°
    sine_table[239] = 16'h9249;  // Angle 239°
    sine_table[240] = 16'h9127;  // Angle 240°
    sine_table[241] = 16'h900D;  // Angle 241°
    sine_table[242] = 16'h8EFC;  // Angle 242°
    sine_table[243] = 16'h8DF4;  // Angle 243°
    sine_table[244] = 16'h8CF5;  // Angle 244°
    sine_table[245] = 16'h8BFF;  // Angle 245°
    sine_table[246] = 16'h8B11;  // Angle 246°
    sine_table[247] = 16'h8A2D;  // Angle 247°
    sine_table[248] = 16'h8953;  // Angle 248°
    sine_table[249] = 16'h8881;  // Angle 249°
    sine_table[250] = 16'h87B9;  // Angle 250°
    sine_table[251] = 16'h86FA;  // Angle 251°
    sine_table[252] = 16'h8644;  // Angle 252°
    sine_table[253] = 16'h8598;  // Angle 253°
    sine_table[254] = 16'h84F6;  // Angle 254°
    sine_table[255] = 16'h845D;  // Angle 255°
    sine_table[256] = 16'h83CE;  // Angle 256°
    sine_table[257] = 16'h8348;  // Angle 257°
    sine_table[258] = 16'h82CD;  // Angle 258°
    sine_table[259] = 16'h825B;  // Angle 259°
    sine_table[260] = 16'h81F2;  // Angle 260°
    sine_table[261] = 16'h8194;  // Angle 261°
    sine_table[262] = 16'h813F;  // Angle 262°
    sine_table[263] = 16'h80F5;  // Angle 263°
    sine_table[264] = 16'h80B4;  // Angle 264°
    sine_table[265] = 16'h807D;  // Angle 265°
    sine_table[266] = 16'h8050;  // Angle 266°
    sine_table[267] = 16'h802D;  // Angle 267°
    sine_table[268] = 16'h8014;  // Angle 268°
    sine_table[269] = 16'h8005;  // Angle 269°
    sine_table[270] = 16'h8000;  // Angle 270°
    sine_table[271] = 16'h8005;  // Angle 271°
    sine_table[272] = 16'h8014;  // Angle 272°
    sine_table[273] = 16'h802D;  // Angle 273°
    sine_table[274] = 16'h8050;  // Angle 274°
    sine_table[275] = 16'h807D;  // Angle 275°
    sine_table[276] = 16'h80B4;  // Angle 276°
    sine_table[277] = 16'h80F5;  // Angle 277°
    sine_table[278] = 16'h813F;  // Angle 278°
    sine_table[279] = 16'h8194;  // Angle 279°
    sine_table[280] = 16'h81F2;  // Angle 280°
    sine_table[281] = 16'h825B;  // Angle 281°
    sine_table[282] = 16'h82CD;  // Angle 282°
    sine_table[283] = 16'h8348;  // Angle 283°
    sine_table[284] = 16'h83CE;  // Angle 284°
    sine_table[285] = 16'h845D;  // Angle 285°
    sine_table[286] = 16'h84F6;  // Angle 286°
    sine_table[287] = 16'h8598;  // Angle 287°
    sine_table[288] = 16'h8644;  // Angle 288°
    sine_table[289] = 16'h86FA;  // Angle 289°
    sine_table[290] = 16'h87B9;  // Angle 290°
    sine_table[291] = 16'h8881;  // Angle 291°
    sine_table[292] = 16'h8953;  // Angle 292°
    sine_table[293] = 16'h8A2D;  // Angle 293°
    sine_table[294] = 16'h8B11;  // Angle 294°
    sine_table[295] = 16'h8BFF;  // Angle 295°
    sine_table[296] = 16'h8CF5;  // Angle 296°
    sine_table[297] = 16'h8DF4;  // Angle 297°
    sine_table[298] = 16'h8EFC;  // Angle 298°
    sine_table[299] = 16'h900D;  // Angle 299°
    sine_table[300] = 16'h9127;  // Angle 300°
    sine_table[301] = 16'h9249;  // Angle 301°
    sine_table[302] = 16'h9374;  // Angle 302°
    sine_table[303] = 16'h94A7;  // Angle 303°
    sine_table[304] = 16'h95E3;  // Angle 304°
    sine_table[305] = 16'h9727;  // Angle 305°
    sine_table[306] = 16'h9873;  // Angle 306°
    sine_table[307] = 16'h99C7;  // Angle 307°
    sine_table[308] = 16'h9B23;  // Angle 308°
    sine_table[309] = 16'h9C87;  // Angle 309°
    sine_table[310] = 16'h9DF3;  // Angle 310°
    sine_table[311] = 16'h9F66;  // Angle 311°
    sine_table[312] = 16'hA0E1;  // Angle 312°
    sine_table[313] = 16'hA264;  // Angle 313°
    sine_table[314] = 16'hA3ED;  // Angle 314°
    sine_table[315] = 16'hA57E;  // Angle 315°
    sine_table[316] = 16'hA716;  // Angle 316°
    sine_table[317] = 16'hA8B5;  // Angle 317°
    sine_table[318] = 16'hAA5A;  // Angle 318°
    sine_table[319] = 16'hAC07;  // Angle 319°
    sine_table[320] = 16'hADBA;  // Angle 320°
    sine_table[321] = 16'hAF73;  // Angle 321°
    sine_table[322] = 16'hB133;  // Angle 322°
    sine_table[323] = 16'hB2F8;  // Angle 323°
    sine_table[324] = 16'hB4C4;  // Angle 324°
    sine_table[325] = 16'hB696;  // Angle 325°
    sine_table[326] = 16'hB86D;  // Angle 326°
    sine_table[327] = 16'hBA4A;  // Angle 327°
    sine_table[328] = 16'hBC2C;  // Angle 328°
    sine_table[329] = 16'hBE14;  // Angle 329°
    sine_table[330] = 16'hC000;  // Angle 330°
    sine_table[331] = 16'hC1F2;  // Angle 331°
    sine_table[332] = 16'hC3E9;  // Angle 332°
    sine_table[333] = 16'hC5E4;  // Angle 333°
    sine_table[334] = 16'hC7E4;  // Angle 334°
    sine_table[335] = 16'hC9E8;  // Angle 335°
    sine_table[336] = 16'hCBF1;  // Angle 336°
    sine_table[337] = 16'hCDFD;  // Angle 337°
    sine_table[338] = 16'hD00D;  // Angle 338°
    sine_table[339] = 16'hD221;  // Angle 339°
    sine_table[340] = 16'hD439;  // Angle 340°
    sine_table[341] = 16'hD654;  // Angle 341°
    sine_table[342] = 16'hD873;  // Angle 342°
    sine_table[343] = 16'hDA94;  // Angle 343°
    sine_table[344] = 16'hDCB8;  // Angle 344°
    sine_table[345] = 16'hDEE0;  // Angle 345°
    sine_table[346] = 16'hE109;  // Angle 346°
    sine_table[347] = 16'hE335;  // Angle 347°
    sine_table[348] = 16'hE564;  // Angle 348°
    sine_table[349] = 16'hE794;  // Angle 349°
    sine_table[350] = 16'hE9C6;  // Angle 350°
    sine_table[351] = 16'hEBFA;  // Angle 351°
    sine_table[352] = 16'hEE30;  // Angle 352°
    sine_table[353] = 16'hF067;  // Angle 353°
    sine_table[354] = 16'hF29F;  // Angle 354°
    sine_table[355] = 16'hF4D9;  // Angle 355°
    sine_table[356] = 16'hF713;  // Angle 356°
    sine_table[357] = 16'hF94E;  // Angle 357°
    sine_table[358] = 16'hFB89;  // Angle 358°
    sine_table[359] = 16'hFDC5;  // Angle 359°

    cosine_table[0] = 16'h7FFF;  // Angle 0°
    cosine_table[1] = 16'h7FFB;  // Angle 1°
    cosine_table[2] = 16'h7FEC;  // Angle 2°
    cosine_table[3] = 16'h7FD3;  // Angle 3°
    cosine_table[4] = 16'h7FB0;  // Angle 4°
    cosine_table[5] = 16'h7F83;  // Angle 5°
    cosine_table[6] = 16'h7F4C;  // Angle 6°
    cosine_table[7] = 16'h7F0B;  // Angle 7°
    cosine_table[8] = 16'h7EC1;  // Angle 8°
    cosine_table[9] = 16'h7E6C;  // Angle 9°
    cosine_table[10] = 16'h7E0E;  // Angle 10°
    cosine_table[11] = 16'h7DA5;  // Angle 11°
    cosine_table[12] = 16'h7D33;  // Angle 12°
    cosine_table[13] = 16'h7CB8;  // Angle 13°
    cosine_table[14] = 16'h7C32;  // Angle 14°
    cosine_table[15] = 16'h7BA3;  // Angle 15°
    cosine_table[16] = 16'h7B0A;  // Angle 16°
    cosine_table[17] = 16'h7A68;  // Angle 17°
    cosine_table[18] = 16'h79BC;  // Angle 18°
    cosine_table[19] = 16'h7906;  // Angle 19°
    cosine_table[20] = 16'h7847;  // Angle 20°
    cosine_table[21] = 16'h777F;  // Angle 21°
    cosine_table[22] = 16'h76AD;  // Angle 22°
    cosine_table[23] = 16'h75D3;  // Angle 23°
    cosine_table[24] = 16'h74EF;  // Angle 24°
    cosine_table[25] = 16'h7401;  // Angle 25°
    cosine_table[26] = 16'h730B;  // Angle 26°
    cosine_table[27] = 16'h720C;  // Angle 27°
    cosine_table[28] = 16'h7104;  // Angle 28°
    cosine_table[29] = 16'h6FF3;  // Angle 29°
    cosine_table[30] = 16'h6ED9;  // Angle 30°
    cosine_table[31] = 16'h6DB7;  // Angle 31°
    cosine_table[32] = 16'h6C8C;  // Angle 32°
    cosine_table[33] = 16'h6B59;  // Angle 33°
    cosine_table[34] = 16'h6A1D;  // Angle 34°
    cosine_table[35] = 16'h68D9;  // Angle 35°
    cosine_table[36] = 16'h678D;  // Angle 36°
    cosine_table[37] = 16'h6639;  // Angle 37°
    cosine_table[38] = 16'h64DD;  // Angle 38°
    cosine_table[39] = 16'h6379;  // Angle 39°
    cosine_table[40] = 16'h620D;  // Angle 40°
    cosine_table[41] = 16'h609A;  // Angle 41°
    cosine_table[42] = 16'h5F1F;  // Angle 42°
    cosine_table[43] = 16'h5D9C;  // Angle 43°
    cosine_table[44] = 16'h5C13;  // Angle 44°
    cosine_table[45] = 16'h5A82;  // Angle 45°
    cosine_table[46] = 16'h58EA;  // Angle 46°
    cosine_table[47] = 16'h574B;  // Angle 47°
    cosine_table[48] = 16'h55A6;  // Angle 48°
    cosine_table[49] = 16'h53F9;  // Angle 49°
    cosine_table[50] = 16'h5246;  // Angle 50°
    cosine_table[51] = 16'h508D;  // Angle 51°
    cosine_table[52] = 16'h4ECD;  // Angle 52°
    cosine_table[53] = 16'h4D08;  // Angle 53°
    cosine_table[54] = 16'h4B3C;  // Angle 54°
    cosine_table[55] = 16'h496A;  // Angle 55°
    cosine_table[56] = 16'h4793;  // Angle 56°
    cosine_table[57] = 16'h45B6;  // Angle 57°
    cosine_table[58] = 16'h43D4;  // Angle 58°
    cosine_table[59] = 16'h41EC;  // Angle 59°
    cosine_table[60] = 16'h4000;  // Angle 60°
    cosine_table[61] = 16'h3E0E;  // Angle 61°
    cosine_table[62] = 16'h3C17;  // Angle 62°
    cosine_table[63] = 16'h3A1C;  // Angle 63°
    cosine_table[64] = 16'h381C;  // Angle 64°
    cosine_table[65] = 16'h3618;  // Angle 65°
    cosine_table[66] = 16'h340F;  // Angle 66°
    cosine_table[67] = 16'h3203;  // Angle 67°
    cosine_table[68] = 16'h2FF3;  // Angle 68°
    cosine_table[69] = 16'h2DDF;  // Angle 69°
    cosine_table[70] = 16'h2BC7;  // Angle 70°
    cosine_table[71] = 16'h29AC;  // Angle 71°
    cosine_table[72] = 16'h278D;  // Angle 72°
    cosine_table[73] = 16'h256C;  // Angle 73°
    cosine_table[74] = 16'h2348;  // Angle 74°
    cosine_table[75] = 16'h2120;  // Angle 75°
    cosine_table[76] = 16'h1EF7;  // Angle 76°
    cosine_table[77] = 16'h1CCB;  // Angle 77°
    cosine_table[78] = 16'h1A9C;  // Angle 78°
    cosine_table[79] = 16'h186C;  // Angle 79°
    cosine_table[80] = 16'h163A;  // Angle 80°
    cosine_table[81] = 16'h1406;  // Angle 81°
    cosine_table[82] = 16'h11D0;  // Angle 82°
    cosine_table[83] = 16'h0F99;  // Angle 83°
    cosine_table[84] = 16'h0D61;  // Angle 84°
    cosine_table[85] = 16'h0B27;  // Angle 85°
    cosine_table[86] = 16'h08ED;  // Angle 86°
    cosine_table[87] = 16'h06B2;  // Angle 87°
    cosine_table[88] = 16'h0477;  // Angle 88°
    cosine_table[89] = 16'h023B;  // Angle 89°
    cosine_table[90] = 16'h0000;  // Angle 90°
    cosine_table[91] = 16'hFDC5;  // Angle 91°
    cosine_table[92] = 16'hFB89;  // Angle 92°
    cosine_table[93] = 16'hF94E;  // Angle 93°
    cosine_table[94] = 16'hF713;  // Angle 94°
    cosine_table[95] = 16'hF4D9;  // Angle 95°
    cosine_table[96] = 16'hF29F;  // Angle 96°
    cosine_table[97] = 16'hF067;  // Angle 97°
    cosine_table[98] = 16'hEE30;  // Angle 98°
    cosine_table[99] = 16'hEBFA;  // Angle 99°
    cosine_table[100] = 16'hE9C6;  // Angle 100°
    cosine_table[101] = 16'hE794;  // Angle 101°
    cosine_table[102] = 16'hE564;  // Angle 102°
    cosine_table[103] = 16'hE335;  // Angle 103°
    cosine_table[104] = 16'hE109;  // Angle 104°
    cosine_table[105] = 16'hDEE0;  // Angle 105°
    cosine_table[106] = 16'hDCB8;  // Angle 106°
    cosine_table[107] = 16'hDA94;  // Angle 107°
    cosine_table[108] = 16'hD873;  // Angle 108°
    cosine_table[109] = 16'hD654;  // Angle 109°
    cosine_table[110] = 16'hD439;  // Angle 110°
    cosine_table[111] = 16'hD221;  // Angle 111°
    cosine_table[112] = 16'hD00D;  // Angle 112°
    cosine_table[113] = 16'hCDFD;  // Angle 113°
    cosine_table[114] = 16'hCBF1;  // Angle 114°
    cosine_table[115] = 16'hC9E8;  // Angle 115°
    cosine_table[116] = 16'hC7E4;  // Angle 116°
    cosine_table[117] = 16'hC5E4;  // Angle 117°
    cosine_table[118] = 16'hC3E9;  // Angle 118°
    cosine_table[119] = 16'hC1F2;  // Angle 119°
    cosine_table[120] = 16'hC001;  // Angle 120°
    cosine_table[121] = 16'hBE14;  // Angle 121°
    cosine_table[122] = 16'hBC2C;  // Angle 122°
    cosine_table[123] = 16'hBA4A;  // Angle 123°
    cosine_table[124] = 16'hB86D;  // Angle 124°
    cosine_table[125] = 16'hB696;  // Angle 125°
    cosine_table[126] = 16'hB4C4;  // Angle 126°
    cosine_table[127] = 16'hB2F8;  // Angle 127°
    cosine_table[128] = 16'hB133;  // Angle 128°
    cosine_table[129] = 16'hAF73;  // Angle 129°
    cosine_table[130] = 16'hADBA;  // Angle 130°
    cosine_table[131] = 16'hAC07;  // Angle 131°
    cosine_table[132] = 16'hAA5A;  // Angle 132°
    cosine_table[133] = 16'hA8B5;  // Angle 133°
    cosine_table[134] = 16'hA716;  // Angle 134°
    cosine_table[135] = 16'hA57E;  // Angle 135°
    cosine_table[136] = 16'hA3ED;  // Angle 136°
    cosine_table[137] = 16'hA264;  // Angle 137°
    cosine_table[138] = 16'hA0E1;  // Angle 138°
    cosine_table[139] = 16'h9F66;  // Angle 139°
    cosine_table[140] = 16'h9DF3;  // Angle 140°
    cosine_table[141] = 16'h9C87;  // Angle 141°
    cosine_table[142] = 16'h9B23;  // Angle 142°
    cosine_table[143] = 16'h99C7;  // Angle 143°
    cosine_table[144] = 16'h9873;  // Angle 144°
    cosine_table[145] = 16'h9727;  // Angle 145°
    cosine_table[146] = 16'h95E3;  // Angle 146°
    cosine_table[147] = 16'h94A7;  // Angle 147°
    cosine_table[148] = 16'h9374;  // Angle 148°
    cosine_table[149] = 16'h9249;  // Angle 149°
    cosine_table[150] = 16'h9127;  // Angle 150°
    cosine_table[151] = 16'h900D;  // Angle 151°
    cosine_table[152] = 16'h8EFC;  // Angle 152°
    cosine_table[153] = 16'h8DF4;  // Angle 153°
    cosine_table[154] = 16'h8CF5;  // Angle 154°
    cosine_table[155] = 16'h8BFF;  // Angle 155°
    cosine_table[156] = 16'h8B11;  // Angle 156°
    cosine_table[157] = 16'h8A2D;  // Angle 157°
    cosine_table[158] = 16'h8953;  // Angle 158°
    cosine_table[159] = 16'h8881;  // Angle 159°
    cosine_table[160] = 16'h87B9;  // Angle 160°
    cosine_table[161] = 16'h86FA;  // Angle 161°
    cosine_table[162] = 16'h8644;  // Angle 162°
    cosine_table[163] = 16'h8598;  // Angle 163°
    cosine_table[164] = 16'h84F6;  // Angle 164°
    cosine_table[165] = 16'h845D;  // Angle 165°
    cosine_table[166] = 16'h83CE;  // Angle 166°
    cosine_table[167] = 16'h8348;  // Angle 167°
    cosine_table[168] = 16'h82CD;  // Angle 168°
    cosine_table[169] = 16'h825B;  // Angle 169°
    cosine_table[170] = 16'h81F2;  // Angle 170°
    cosine_table[171] = 16'h8194;  // Angle 171°
    cosine_table[172] = 16'h813F;  // Angle 172°
    cosine_table[173] = 16'h80F5;  // Angle 173°
    cosine_table[174] = 16'h80B4;  // Angle 174°
    cosine_table[175] = 16'h807D;  // Angle 175°
    cosine_table[176] = 16'h8050;  // Angle 176°
    cosine_table[177] = 16'h802D;  // Angle 177°
    cosine_table[178] = 16'h8014;  // Angle 178°
    cosine_table[179] = 16'h8005;  // Angle 179°
    cosine_table[180] = 16'h8000;  // Angle 180°
    cosine_table[181] = 16'h8005;  // Angle 181°
    cosine_table[182] = 16'h8014;  // Angle 182°
    cosine_table[183] = 16'h802D;  // Angle 183°
    cosine_table[184] = 16'h8050;  // Angle 184°
    cosine_table[185] = 16'h807D;  // Angle 185°
    cosine_table[186] = 16'h80B4;  // Angle 186°
    cosine_table[187] = 16'h80F5;  // Angle 187°
    cosine_table[188] = 16'h813F;  // Angle 188°
    cosine_table[189] = 16'h8194;  // Angle 189°
    cosine_table[190] = 16'h81F2;  // Angle 190°
    cosine_table[191] = 16'h825B;  // Angle 191°
    cosine_table[192] = 16'h82CD;  // Angle 192°
    cosine_table[193] = 16'h8348;  // Angle 193°
    cosine_table[194] = 16'h83CE;  // Angle 194°
    cosine_table[195] = 16'h845D;  // Angle 195°
    cosine_table[196] = 16'h84F6;  // Angle 196°
    cosine_table[197] = 16'h8598;  // Angle 197°
    cosine_table[198] = 16'h8644;  // Angle 198°
    cosine_table[199] = 16'h86FA;  // Angle 199°
    cosine_table[200] = 16'h87B9;  // Angle 200°
    cosine_table[201] = 16'h8881;  // Angle 201°
    cosine_table[202] = 16'h8953;  // Angle 202°
    cosine_table[203] = 16'h8A2D;  // Angle 203°
    cosine_table[204] = 16'h8B11;  // Angle 204°
    cosine_table[205] = 16'h8BFF;  // Angle 205°
    cosine_table[206] = 16'h8CF5;  // Angle 206°
    cosine_table[207] = 16'h8DF4;  // Angle 207°
    cosine_table[208] = 16'h8EFC;  // Angle 208°
    cosine_table[209] = 16'h900D;  // Angle 209°
    cosine_table[210] = 16'h9127;  // Angle 210°
    cosine_table[211] = 16'h9249;  // Angle 211°
    cosine_table[212] = 16'h9374;  // Angle 212°
    cosine_table[213] = 16'h94A7;  // Angle 213°
    cosine_table[214] = 16'h95E3;  // Angle 214°
    cosine_table[215] = 16'h9727;  // Angle 215°
    cosine_table[216] = 16'h9873;  // Angle 216°
    cosine_table[217] = 16'h99C7;  // Angle 217°
    cosine_table[218] = 16'h9B23;  // Angle 218°
    cosine_table[219] = 16'h9C87;  // Angle 219°
    cosine_table[220] = 16'h9DF3;  // Angle 220°
    cosine_table[221] = 16'h9F66;  // Angle 221°
    cosine_table[222] = 16'hA0E1;  // Angle 222°
    cosine_table[223] = 16'hA264;  // Angle 223°
    cosine_table[224] = 16'hA3ED;  // Angle 224°
    cosine_table[225] = 16'hA57E;  // Angle 225°
    cosine_table[226] = 16'hA716;  // Angle 226°
    cosine_table[227] = 16'hA8B5;  // Angle 227°
    cosine_table[228] = 16'hAA5A;  // Angle 228°
    cosine_table[229] = 16'hAC07;  // Angle 229°
    cosine_table[230] = 16'hADBA;  // Angle 230°
    cosine_table[231] = 16'hAF73;  // Angle 231°
    cosine_table[232] = 16'hB133;  // Angle 232°
    cosine_table[233] = 16'hB2F8;  // Angle 233°
    cosine_table[234] = 16'hB4C4;  // Angle 234°
    cosine_table[235] = 16'hB696;  // Angle 235°
    cosine_table[236] = 16'hB86D;  // Angle 236°
    cosine_table[237] = 16'hBA4A;  // Angle 237°
    cosine_table[238] = 16'hBC2C;  // Angle 238°
    cosine_table[239] = 16'hBE14;  // Angle 239°
    cosine_table[240] = 16'hC000;  // Angle 240°
    cosine_table[241] = 16'hC1F2;  // Angle 241°
    cosine_table[242] = 16'hC3E9;  // Angle 242°
    cosine_table[243] = 16'hC5E4;  // Angle 243°
    cosine_table[244] = 16'hC7E4;  // Angle 244°
    cosine_table[245] = 16'hC9E8;  // Angle 245°
    cosine_table[246] = 16'hCBF1;  // Angle 246°
    cosine_table[247] = 16'hCDFD;  // Angle 247°
    cosine_table[248] = 16'hD00D;  // Angle 248°
    cosine_table[249] = 16'hD221;  // Angle 249°
    cosine_table[250] = 16'hD439;  // Angle 250°
    cosine_table[251] = 16'hD654;  // Angle 251°
    cosine_table[252] = 16'hD873;  // Angle 252°
    cosine_table[253] = 16'hDA94;  // Angle 253°
    cosine_table[254] = 16'hDCB8;  // Angle 254°
    cosine_table[255] = 16'hDEE0;  // Angle 255°
    cosine_table[256] = 16'hE109;  // Angle 256°
    cosine_table[257] = 16'hE335;  // Angle 257°
    cosine_table[258] = 16'hE564;  // Angle 258°
    cosine_table[259] = 16'hE794;  // Angle 259°
    cosine_table[260] = 16'hE9C6;  // Angle 260°
    cosine_table[261] = 16'hEBFA;  // Angle 261°
    cosine_table[262] = 16'hEE30;  // Angle 262°
    cosine_table[263] = 16'hF067;  // Angle 263°
    cosine_table[264] = 16'hF29F;  // Angle 264°
    cosine_table[265] = 16'hF4D9;  // Angle 265°
    cosine_table[266] = 16'hF713;  // Angle 266°
    cosine_table[267] = 16'hF94E;  // Angle 267°
    cosine_table[268] = 16'hFB89;  // Angle 268°
    cosine_table[269] = 16'hFDC5;  // Angle 269°
    cosine_table[270] = 16'h0000;  // Angle 270°
    cosine_table[271] = 16'h023B;  // Angle 271°
    cosine_table[272] = 16'h0477;  // Angle 272°
    cosine_table[273] = 16'h06B2;  // Angle 273°
    cosine_table[274] = 16'h08ED;  // Angle 274°
    cosine_table[275] = 16'h0B27;  // Angle 275°
    cosine_table[276] = 16'h0D61;  // Angle 276°
    cosine_table[277] = 16'h0F99;  // Angle 277°
    cosine_table[278] = 16'h11D0;  // Angle 278°
    cosine_table[279] = 16'h1406;  // Angle 279°
    cosine_table[280] = 16'h163A;  // Angle 280°
    cosine_table[281] = 16'h186C;  // Angle 281°
    cosine_table[282] = 16'h1A9C;  // Angle 282°
    cosine_table[283] = 16'h1CCB;  // Angle 283°
    cosine_table[284] = 16'h1EF7;  // Angle 284°
    cosine_table[285] = 16'h2120;  // Angle 285°
    cosine_table[286] = 16'h2348;  // Angle 286°
    cosine_table[287] = 16'h256C;  // Angle 287°
    cosine_table[288] = 16'h278D;  // Angle 288°
    cosine_table[289] = 16'h29AC;  // Angle 289°
    cosine_table[290] = 16'h2BC7;  // Angle 290°
    cosine_table[291] = 16'h2DDF;  // Angle 291°
    cosine_table[292] = 16'h2FF3;  // Angle 292°
    cosine_table[293] = 16'h3203;  // Angle 293°
    cosine_table[294] = 16'h340F;  // Angle 294°
    cosine_table[295] = 16'h3618;  // Angle 295°
    cosine_table[296] = 16'h381C;  // Angle 296°
    cosine_table[297] = 16'h3A1C;  // Angle 297°
    cosine_table[298] = 16'h3C17;  // Angle 298°
    cosine_table[299] = 16'h3E0E;  // Angle 299°
    cosine_table[300] = 16'h4000;  // Angle 300°
    cosine_table[301] = 16'h41EC;  // Angle 301°
    cosine_table[302] = 16'h43D4;  // Angle 302°
    cosine_table[303] = 16'h45B6;  // Angle 303°
    cosine_table[304] = 16'h4793;  // Angle 304°
    cosine_table[305] = 16'h496A;  // Angle 305°
    cosine_table[306] = 16'h4B3C;  // Angle 306°
    cosine_table[307] = 16'h4D08;  // Angle 307°
    cosine_table[308] = 16'h4ECD;  // Angle 308°
    cosine_table[309] = 16'h508D;  // Angle 309°
    cosine_table[310] = 16'h5246;  // Angle 310°
    cosine_table[311] = 16'h53F9;  // Angle 311°
    cosine_table[312] = 16'h55A6;  // Angle 312°
    cosine_table[313] = 16'h574B;  // Angle 313°
    cosine_table[314] = 16'h58EA;  // Angle 314°
    cosine_table[315] = 16'h5A82;  // Angle 315°
    cosine_table[316] = 16'h5C13;  // Angle 316°
    cosine_table[317] = 16'h5D9C;  // Angle 317°
    cosine_table[318] = 16'h5F1F;  // Angle 318°
    cosine_table[319] = 16'h609A;  // Angle 319°
    cosine_table[320] = 16'h620D;  // Angle 320°
    cosine_table[321] = 16'h6379;  // Angle 321°
    cosine_table[322] = 16'h64DD;  // Angle 322°
    cosine_table[323] = 16'h6639;  // Angle 323°
    cosine_table[324] = 16'h678D;  // Angle 324°
    cosine_table[325] = 16'h68D9;  // Angle 325°
    cosine_table[326] = 16'h6A1D;  // Angle 326°
    cosine_table[327] = 16'h6B59;  // Angle 327°
    cosine_table[328] = 16'h6C8C;  // Angle 328°
    cosine_table[329] = 16'h6DB7;  // Angle 329°
    cosine_table[330] = 16'h6ED9;  // Angle 330°
    cosine_table[331] = 16'h6FF3;  // Angle 331°
    cosine_table[332] = 16'h7104;  // Angle 332°
    cosine_table[333] = 16'h720C;  // Angle 333°
    cosine_table[334] = 16'h730B;  // Angle 334°
    cosine_table[335] = 16'h7401;  // Angle 335°
    cosine_table[336] = 16'h74EF;  // Angle 336°
    cosine_table[337] = 16'h75D3;  // Angle 337°
    cosine_table[338] = 16'h76AD;  // Angle 338°
    cosine_table[339] = 16'h777F;  // Angle 339°
    cosine_table[340] = 16'h7847;  // Angle 340°
    cosine_table[341] = 16'h7906;  // Angle 341°
    cosine_table[342] = 16'h79BC;  // Angle 342°
    cosine_table[343] = 16'h7A68;  // Angle 343°
    cosine_table[344] = 16'h7B0A;  // Angle 344°
    cosine_table[345] = 16'h7BA3;  // Angle 345°
    cosine_table[346] = 16'h7C32;  // Angle 346°
    cosine_table[347] = 16'h7CB8;  // Angle 347°
    cosine_table[348] = 16'h7D33;  // Angle 348°
    cosine_table[349] = 16'h7DA5;  // Angle 349°
    cosine_table[350] = 16'h7E0E;  // Angle 350°
    cosine_table[351] = 16'h7E6C;  // Angle 351°
    cosine_table[352] = 16'h7EC1;  // Angle 352°
    cosine_table[353] = 16'h7F0B;  // Angle 353°
    cosine_table[354] = 16'h7F4C;  // Angle 354°
    cosine_table[355] = 16'h7F83;  // Angle 355°
    cosine_table[356] = 16'h7FB0;  // Angle 356°
    cosine_table[357] = 16'h7FD3;  // Angle 357°
    cosine_table[358] = 16'h7FEC;  // Angle 358°
    cosine_table[359] = 16'h7FFB;  // Angle 359°
  end

  // Output sine and cosine based on the angle
  always @(*) begin
    sine_out = sine_table[angle];
    cosine_out = cosine_table[angle];
  end

endmodule
