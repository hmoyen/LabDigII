// module angle_to_coordinates(
//     input [6:0] angle,  // 7-bit input (0 to 90 degrees)
//     output reg [16:0] x,
//     output reg [16:0] y,
//     output reg [16:0] z
// );

//     // ROM for coordinates
//     reg [16:0] x_rom [0:127];
//     reg [16:0] y_rom [0:127];
//     reg [16:0] z_rom [0:127];

//     initial begin
//         // Initializ_rome the ROM with the given values (only_rom a portion shown for brevity_rom)
//         x_rom[0] <= 17'd32768;  y_rom[0] <= 17'd0;      z_rom[0] <= 17'd0;
//         x_rom[1] <= 17'd32763;  y_rom[1] <= 17'd571;    z_rom[1] <= 17'd571;
//         x_rom[2] <= 17'd32748;  y_rom[2] <= 17'd1143;   z_rom[2] <= 17'd1143;
//         x_rom[3] <= 17'd32723;  y_rom[3] <= 17'd1714;   z_rom[3] <= 17'd1715;
//         x_rom[4] <= 17'd32688;  y_rom[4] <= 17'd2285;   z_rom[4] <= 17'd2287;
//         x_rom[5] <= 17'd32643;  y_rom[5] <= 17'd2855;   z_rom[5] <= 17'd2859;
//         x_rom[6] <= 17'd32588;  y_rom[6] <= 17'd3425;   z_rom[6] <= 17'd3431;
//         x_rom[7] <= 17'd32523;  y_rom[7] <= 17'd3993;   z_rom[7] <= 17'd4003;
//         x_rom[8] <= 17'd32449;  y_rom[8] <= 17'd4560;   z_rom[8] <= 17'd4575;
//         x_rom[9] <= 17'd32364;  y_rom[9] <= 17'd5126;   z_rom[9] <= 17'd5147;
//         x_rom[10] <= 17'd32270; y_rom[10] <= 17'd5690;  z_rom[10] <= 17'd5719;
//         x_rom[11] <= 17'd32165; y_rom[11] <= 17'd6252;  z_rom[11] <= 17'd6291;
//         x_rom[12] <= 17'd32051; y_rom[12] <= 17'd6812;  z_rom[12] <= 17'd6862;
//         x_rom[13] <= 17'd31928; y_rom[13] <= 17'd7371;  z_rom[13] <= 17'd7434;
//         x_rom[14] <= 17'd31794; y_rom[14] <= 17'd7927;  z_rom[14] <= 17'd8006;
//         x_rom[15] <= 17'd31651; y_rom[15] <= 17'd8480;  z_rom[15] <= 17'd8578;
//         x_rom[16] <= 17'd31498; y_rom[16] <= 17'd9032;  z_rom[16] <= 17'd9150;
//         x_rom[17] <= 17'd31336; y_rom[17] <= 17'd9580;  z_rom[17] <= 17'd9722;
//         x_rom[18] <= 17'd31164; y_rom[18] <= 17'd10125; z_rom[18] <= 17'd10294;
//         x_rom[19] <= 17'd30982; y_rom[19] <= 17'd10668; z_rom[19] <= 17'd10866;
//         x_rom[20] <= 17'd30791; y_rom[20] <= 17'd11207; z_rom[20] <= 17'd11438;
//         x_rom[21] <= 17'd30591; y_rom[21] <= 17'd11743; z_rom[21] <= 17'd12010;
//         x_rom[22] <= 17'd30381; y_rom[22] <= 17'd12275; z_rom[22] <= 17'd12582;
//         x_rom[23] <= 17'd30163; y_rom[23] <= 17'd12803; z_rom[23] <= 17'd13153;
//         x_rom[24] <= 17'd29935; y_rom[24] <= 17'd13327; z_rom[24] <= 17'd13725;
//         x_rom[25] <= 17'd29697; y_rom[25] <= 17'd13848; z_rom[25] <= 17'd14297;
//         x_rom[26] <= 17'd29451; y_rom[26] <= 17'd14364; z_rom[26] <= 17'd14869;
//         x_rom[27] <= 17'd29196; y_rom[27] <= 17'd14876; z_rom[27] <= 17'd15441;
//         x_rom[28] <= 17'd28932; y_rom[28] <= 17'd15383; z_rom[28] <= 17'd16013;
//         x_rom[29] <= 17'd28659; y_rom[29] <= 17'd15886; z_rom[29] <= 17'd16585;
//         x_rom[30] <= 17'd28377; y_rom[30] <= 17'd16383; z_rom[30] <= 17'd17157;
//         x_rom[31] <= 17'd28087; y_rom[31] <= 17'd16876; z_rom[31] <= 17'd17729;
//         x_rom[32] <= 17'd27788; y_rom[32] <= 17'd17364; z_rom[32] <= 17'd18301;
//         x_rom[33] <= 17'd27481; y_rom[33] <= 17'd17846; z_rom[33] <= 17'd18873;
//         x_rom[34] <= 17'd27165; y_rom[34] <= 17'd18323; z_rom[34] <= 17'd19444;
//         x_rom[35] <= 17'd26841; y_rom[35] <= 17'd18794; z_rom[35] <= 17'd20016;
//         x_rom[36] <= 17'd26509; y_rom[36] <= 17'd19260; z_rom[36] <= 17'd20588;
//         x_rom[37] <= 17'd26169; y_rom[37] <= 17'd19720; z_rom[37] <= 17'd21160;
//         x_rom[38] <= 17'd25821; y_rom[38] <= 17'd20173; z_rom[38] <= 17'd21732;
//         x_rom[39] <= 17'd25465; y_rom[39] <= 17'd20621; z_rom[39] <= 17'd22304;
//         x_rom[40] <= 17'd25101; y_rom[40] <= 17'd21062; z_rom[40] <= 17'd22876;
//         x_rom[41] <= 17'd24730; y_rom[41] <= 17'd21497; z_rom[41] <= 17'd23448;
//         x_rom[42] <= 17'd24351; y_rom[42] <= 17'd21926; z_rom[42] <= 17'd24020;
//         x_rom[43] <= 17'd23964; y_rom[43] <= 17'd22347; z_rom[43] <= 17'd24592;
//         x_rom[44] <= 17'd23571; y_rom[44] <= 17'd22762; z_rom[44] <= 17'd25164;
//         x_rom[45] <= 17'd23170; y_rom[45] <= 17'd23170; z_rom[45] <= 17'd25735;
//         x_rom[46] <= 17'd22762; y_rom[46] <= 17'd23571; z_rom[46] <= 17'd26307;
//         x_rom[47] <= 17'd22347; y_rom[47] <= 17'd23964; z_rom[47] <= 17'd26879;
//         x_rom[48] <= 17'd21926; y_rom[48] <= 17'd24351; z_rom[48] <= 17'd27451;
//         x_rom[49] <= 17'd21497; y_rom[49] <= 17'd24730; z_rom[49] <= 17'd28023;
//         x_rom[50] <= 17'd21062; y_rom[50] <= 17'd25101; z_rom[50] <= 17'd28595;
//         x_rom[51] <= 17'd20621; y_rom[51] <= 17'd25465; z_rom[51] <= 17'd29167;
//         x_rom[52] <= 17'd20173; y_rom[52] <= 17'd25821; z_rom[52] <= 17'd29739;
//         x_rom[53] <= 17'd19720; y_rom[53] <= 17'd26169; z_rom[53] <= 17'd30311;
//         x_rom[54] <= 17'd19260; y_rom[54] <= 17'd26509; z_rom[54] <= 17'd30883;
//         x_rom[55] <= 17'd18794; y_rom[55] <= 17'd26841; z_rom[55] <= 17'd31455;
//         x_rom[56] <= 17'd18323; y_rom[56] <= 17'd27165; z_rom[56] <= 17'd32026;
//         x_rom[57] <= 17'd17846; y_rom[57] <= 17'd27481; z_rom[57] <= 17'd32598;
//         x_rom[58] <= 17'd17364; y_rom[58] <= 17'd27788; z_rom[58] <= 17'd33170;
//         x_rom[59] <= 17'd16876; y_rom[59] <= 17'd28087; z_rom[59] <= 17'd33742;
//         x_rom[60] <= 17'd16384; y_rom[60] <= 17'd28377; z_rom[60] <= 17'd34314;
//         x_rom[61] <= 17'd15886; y_rom[61] <= 17'd28659; z_rom[61] <= 17'd34886;
//         x_rom[62] <= 17'd15383; y_rom[62] <= 17'd28932; z_rom[62] <= 17'd35458;
//         x_rom[63] <= 17'd14876; y_rom[63] <= 17'd29196; z_rom[63] <= 17'd36030;
//         x_rom[64] <= 17'd14364; y_rom[64] <= 17'd29451; z_rom[64] <= 17'd36602;
//         x_rom[65] <= 17'd13848; y_rom[65] <= 17'd29697; z_rom[65] <= 17'd37174;
//         x_rom[66] <= 17'd13327; y_rom[66] <= 17'd29935; z_rom[66] <= 17'd37746;
//         x_rom[67] <= 17'd12803; y_rom[67] <= 17'd30163; z_rom[67] <= 17'd38317;
//         x_rom[68] <= 17'd12275; y_rom[68] <= 17'd30381; z_rom[68] <= 17'd38889;
//         x_rom[69] <= 17'd11743; y_rom[69] <= 17'd30591; z_rom[69] <= 17'd39461;
//         x_rom[70] <= 17'd11207; y_rom[70] <= 17'd30791; z_rom[70] <= 17'd40033;
//         x_rom[71] <= 17'd10668; y_rom[71] <= 17'd30982; z_rom[71] <= 17'd40605;
//         x_rom[72] <= 17'd10125; y_rom[72] <= 17'd31164; z_rom[72] <= 17'd41177;
//         x_rom[73] <= 17'd9580;  y_rom[73] <= 17'd31336; z_rom[73] <= 17'd41749;
//         x_rom[74] <= 17'd9032;  y_rom[74] <= 17'd31498; z_rom[74] <= 17'd42321;
//         x_rom[75] <= 17'd8480;  y_rom[75] <= 17'd31651; z_rom[75] <= 17'd42893;
//         x_rom[76] <= 17'd7927;  y_rom[76] <= 17'd31794; z_rom[76] <= 17'd43465;
//         x_rom[77] <= 17'd7371;  y_rom[77] <= 17'd31928; z_rom[77] <= 17'd44037;
//         x_rom[78] <= 17'd6812;  y_rom[78] <= 17'd32051; z_rom[78] <= 17'd44608;
//         x_rom[79] <= 17'd6252;  y_rom[79] <= 17'd32165; z_rom[79] <= 17'd45180;
//         x_rom[80] <= 17'd5690;  y_rom[80] <= 17'd32270; z_rom[80] <= 17'd45752;
//         x_rom[81] <= 17'd5126;  y_rom[81] <= 17'd32364; z_rom[81] <= 17'd46324;
//         x_rom[82] <= 17'd4560;  y_rom[82] <= 17'd32449; z_rom[82] <= 17'd46896;
//         x_rom[83] <= 17'd3993;  y_rom[83] <= 17'd32523; z_rom[83] <= 17'd47468;
//         x_rom[84] <= 17'd3425;  y_rom[84] <= 17'd32588; z_rom[84] <= 17'd48040;
//         x_rom[85] <= 17'd2855;  y_rom[85] <= 17'd32643; z_rom[85] <= 17'd48612;
//         x_rom[86] <= 17'd2285;  y_rom[86] <= 17'd32688; z_rom[86] <= 17'd49184;
//         x_rom[87] <= 17'd1714;  y_rom[87] <= 17'd32723; z_rom[87] <= 17'd49756;
//         x_rom[88] <= 17'd1143;  y_rom[88] <= 17'd32748; z_rom[88] <= 17'd50328;
//         x_rom[89] <= 17'd571;   y_rom[89] <= 17'd32763; z_rom[89] <= 17'd50899;
//         x_rom[90] <= 17'd0;     y_rom[90] <= 17'd32768; z_rom[90] <= 17'd51471;
//     end

//     alway_roms @(*) begin
//         if (angle <= 90) begin
//             x_rom = x_rom_rom[angle];
//             y_rom = y_rom_rom[angle];
//             z_rom = z_rom_rom[angle];
//         end else begin
//             x_rom = 17'd0;
//             y_rom = 17'd0;
//             z_rom = 17'd0;  // Default value for out of range
//         end
//     end
// endmodule
